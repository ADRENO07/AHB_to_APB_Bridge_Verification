class ahb_master_sequencer extends uvm_sequencer#(ahb_mxtn);
	`uvm_component_utils(ahb_master_sequencer)

	function new(string name = "ahb_master_sequencer", uvm_component parent);
		super.new(name,parent);
	endfunction
endclass
